module aes_encryptor_block();

endmodule 