module AES_Decryptor();
endmodule 